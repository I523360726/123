//============================================================
//Module   : symbol measure
//Function : measure symbol len
//File Tree: 
//-------------------------------------------------------------
//Update History
//-------------------------------------------------------------
//Rev.level     Date          Code_by         Contents
//1.0           2022/11/6     xxxx            Create
//=============================================================
module symbol_measure #(
    `include "com_param.svh"
    parameter END_OF_LIST = 1
)(

);
  
endmodule
